library verilog;
use verilog.vl_types.all;
entity component_test_vlg_vec_tst is
end component_test_vlg_vec_tst;
